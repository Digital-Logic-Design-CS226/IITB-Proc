library work;
use work.all;


library IEEE;
use ieee.std_logic_1164.all;

entity Testbench1 is
end Testbench1;

architecture tb of Testbench1 is
	signal clk, rst: std_logic;
	signal reg_0, reg_1, reg_2, reg_3, reg_4, reg_5, reg_6, reg_7 : std_logic_vector(15 downto 0);
	signal PC_out_1 : std_logic_vector(15 downto 0);
	signal Instruction_returned : std_logic_vector(15 downto 0);
	signal cpc_wrt, cir_write , creg_read,  creg_write,  cpc_update ,  cstatus_reg_write, cLA_SA_reg_write , cmem_read , cmem_write : std_logic;
	signal cwhich_reg : std_logic_vector(2 downto 0);
	signal cSA_which_reg_control : std_logic;
	signal opcode_out : std_logic_vector(3 downto 0);
	signal indata_received : std_logic_vector (15 downto 0);
	signal data_RF_out : std_logic_vector(15 downto 0);
	signal ALU_output_tb : std_logic_vector(15 downto 0);
	signal ALU_A_out : std_logic_vector (15 downto 0);
	signal ALU_B_out : std_logic_vector (15 downto 0);	

	
	component RISC is
	port ( rst: in std_logic;
	indata_received : out std_logic_vector (15 downto 0);
reg_0 : out std_logic_vector(15 downto 0);
reg_1 : out std_logic_vector(15 downto 0);
reg_2 : out std_logic_vector(15 downto 0);
reg_3 : out std_logic_vector(15 downto 0);
reg_4 : out std_logic_vector(15 downto 0);
reg_5 : out std_logic_vector(15 downto 0);
reg_6 : out std_logic_vector(15 downto 0);
reg_7 : out std_logic_vector(15 downto 0);
PC_out_1 : out std_logic_vector(15 downto 0);
Instruction_returned : out std_logic_vector(15 downto 0);
cpc_wrt : out std_logic;
cir_write : out std_logic;
creg_read : out std_logic;
creg_write : out std_logic;
cpc_update : out std_logic;
cstatus_reg_write : out std_logic;
cLA_SA_reg_write : out std_logic;
cmem_read : out std_logic;
cmem_write : out std_logic;
cwhich_reg : out std_logic_vector(2 downto 0);
cSA_which_reg_control : out std_logic;
opcode_out : out std_logic_vector(3 downto 0);
data_RF_out : out std_logic_vector(15 downto 0);
ALU_output_tb : out std_logic_vector(15 downto 0);
ALU_A_out : out std_logic_vector (15 downto 0);
ALU_B_out : out std_logic_vector (15 downto 0);
clk: in std_logic);

	end component;

	begin
	dut_instance: RISC
--	port map(rst, clk);
	port map(rst => rst, indata_received => indata_received, reg_0 => reg_0, reg_1 => reg_1, reg_2 => reg_2, reg_3 => reg_3, reg_4 => reg_4, reg_5 => reg_5, reg_6 => reg_6, reg_7 => reg_7, PC_out_1 => PC_out_1, Instruction_returned => Instruction_returned,  
	cpc_wrt => cpc_wrt, cir_write => cir_write , creg_read => creg_read,  creg_write => creg_write,  cpc_update => cpc_update ,  cstatus_reg_write => cstatus_reg_write, cLA_SA_reg_write => cLA_SA_reg_write , cmem_read => cmem_read , cmem_write => cmem_write,
	cwhich_reg => cwhich_reg,
	cSA_which_reg_control => cSA_which_reg_control,	opcode_out => opcode_out, data_RF_out => data_RF_out, ALU_output_tb => ALU_output_tb,
	ALU_A_out => ALU_A_out, ALU_B_out => ALU_B_out, clk => clk);
	process
	begin
	
	clk<='0';
	rst<='1';
	wait for 10 ns;
	clk<='1';
	rst<='1';
	wait for 10 ns;
	
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	
	
	end process;
end tb;