library work;
use work.all;


library IEEE;
use ieee.std_logic_1164.all;

entity Testbench1 is
end Testbench1;

architecture tb of Testbench1 is
	signal clk, rst: std_logic;
	
	component RISC is
	port ( clk, rst : in std_logic );
	end component;

	begin
	dut_instance: RST
	port map(clk => clk, rst => rst);
	process
	begin
	
	clk<='0';
	rst<='1';
	wait for 10 ns;
	clk<='1';
	rst<='1';
	wait for 10 ns;
	
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	 clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	clk<='0';
	rst<='0';
	wait for 10 ns;
	clk<='1';
	rst<='0';
	wait for 10 ns;
	
	
	end process;
end tb;